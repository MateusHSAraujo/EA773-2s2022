library verilog;
use verilog.vl_types.all;
entity rom16x8_00_vlg_vec_tst is
end rom16x8_00_vlg_vec_tst;
