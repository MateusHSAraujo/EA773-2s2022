library verilog;
use verilog.vl_types.all;
entity bus_tristate_vlg_vec_tst is
end bus_tristate_vlg_vec_tst;
