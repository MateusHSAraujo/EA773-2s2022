library verilog;
use verilog.vl_types.all;
entity computador_simplificado_vlg_vec_tst is
end computador_simplificado_vlg_vec_tst;
