library verilog;
use verilog.vl_types.all;
entity somador_4_bits_vlg_vec_tst is
end somador_4_bits_vlg_vec_tst;
