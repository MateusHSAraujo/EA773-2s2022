library verilog;
use verilog.vl_types.all;
entity rom64x8_0_vlg_vec_tst is
end rom64x8_0_vlg_vec_tst;
