library verilog;
use verilog.vl_types.all;
entity Testemux8x4_vlg_vec_tst is
end Testemux8x4_vlg_vec_tst;
