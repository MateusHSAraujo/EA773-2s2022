library verilog;
use verilog.vl_types.all;
entity decoderBIN_ONEH_vlg_vec_tst is
end decoderBIN_ONEH_vlg_vec_tst;
