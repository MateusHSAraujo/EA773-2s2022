library verilog;
use verilog.vl_types.all;
entity rom16x4_0_vlg_vec_tst is
end rom16x4_0_vlg_vec_tst;
