library verilog;
use verilog.vl_types.all;
entity meio_somador_vlg_sample_tst is
    port(
        xi              : in     vl_logic;
        yi              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end meio_somador_vlg_sample_tst;
