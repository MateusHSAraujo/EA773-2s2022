library verilog;
use verilog.vl_types.all;
entity bus_decodificador_7seg_vlg_vec_tst is
end bus_decodificador_7seg_vlg_vec_tst;
