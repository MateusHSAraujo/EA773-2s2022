library verilog;
use verilog.vl_types.all;
entity bus_ula_vlg_vec_tst is
end bus_ula_vlg_vec_tst;
