library verilog;
use verilog.vl_types.all;
entity rom16x4_2ls_vlg_vec_tst is
end rom16x4_2ls_vlg_vec_tst;
