library verilog;
use verilog.vl_types.all;
entity projeto2_vlg_vec_tst is
end projeto2_vlg_vec_tst;
