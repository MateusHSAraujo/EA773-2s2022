library verilog;
use verilog.vl_types.all;
entity contador_mod_256_vlg_vec_tst is
end contador_mod_256_vlg_vec_tst;
