library verilog;
use verilog.vl_types.all;
entity memprog_vlg_check_tst is
    port(
        drom            : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end memprog_vlg_check_tst;
