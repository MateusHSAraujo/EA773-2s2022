library verilog;
use verilog.vl_types.all;
entity rom64x8_3_vlg_vec_tst is
end rom64x8_3_vlg_vec_tst;
