library verilog;
use verilog.vl_types.all;
entity ram1x4_vlg_vec_tst is
end ram1x4_vlg_vec_tst;
