library verilog;
use verilog.vl_types.all;
entity rom32x8_par10101010impar01010101_vlg_vec_tst is
end rom32x8_par10101010impar01010101_vlg_vec_tst;
