library verilog;
use verilog.vl_types.all;
entity registrador_4_bits_vlg_vec_tst is
end registrador_4_bits_vlg_vec_tst;
