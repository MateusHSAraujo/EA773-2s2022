library verilog;
use verilog.vl_types.all;
entity memprog_vlg_vec_tst is
end memprog_vlg_vec_tst;
