library verilog;
use verilog.vl_types.all;
entity mux16x4_vlg_vec_tst is
end mux16x4_vlg_vec_tst;
