library verilog;
use verilog.vl_types.all;
entity decod_inst_trf_interno_vlg_vec_tst is
end decod_inst_trf_interno_vlg_vec_tst;
