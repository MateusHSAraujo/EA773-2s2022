library verilog;
use verilog.vl_types.all;
entity Testemux16x8_vlg_vec_tst is
end Testemux16x8_vlg_vec_tst;
