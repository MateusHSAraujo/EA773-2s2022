library verilog;
use verilog.vl_types.all;
entity rom32x8_2_vlg_vec_tst is
end rom32x8_2_vlg_vec_tst;
