library verilog;
use verilog.vl_types.all;
entity rom_4blocks_vlg_vec_tst is
end rom_4blocks_vlg_vec_tst;
