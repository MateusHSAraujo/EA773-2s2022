library verilog;
use verilog.vl_types.all;
entity projeto1_vlg_vec_tst is
end projeto1_vlg_vec_tst;
