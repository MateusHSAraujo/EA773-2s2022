library verilog;
use verilog.vl_types.all;
entity meio_somador_vlg_check_tst is
    port(
        gi              : in     vl_logic;
        pi              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end meio_somador_vlg_check_tst;
