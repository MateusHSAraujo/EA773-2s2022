library verilog;
use verilog.vl_types.all;
entity decod_inst_art_vlg_vec_tst is
end decod_inst_art_vlg_vec_tst;
