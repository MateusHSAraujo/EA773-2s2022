library verilog;
use verilog.vl_types.all;
entity rom16x8_zerada_vlg_vec_tst is
end rom16x8_zerada_vlg_vec_tst;
