library verilog;
use verilog.vl_types.all;
entity teste_RAM_vlg_sample_tst is
    port(
        KEY             : in     vl_logic_vector(0 downto 0);
        sampler_tx      : out    vl_logic
    );
end teste_RAM_vlg_sample_tst;
