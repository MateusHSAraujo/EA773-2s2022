library verilog;
use verilog.vl_types.all;
entity somador_completo_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        zi              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end somador_completo_vlg_check_tst;
