library verilog;
use verilog.vl_types.all;
entity Testemux16x4_vlg_vec_tst is
end Testemux16x4_vlg_vec_tst;
